library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use ieee.numeric_std.all;

entity CTRL is
	port(	
		clk_25	: in std_logic;
		CLK		: out std_logic;
		D0			: out std_logic;
		D1			: out std_logic;
		D2			: out std_logic
	);
end entity;


architecture struct of CTRL is


begin
	
		
end;









